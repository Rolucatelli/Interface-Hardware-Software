
module memoria(pc, out);

    input [5:0] pc;
    output reg [15:0] out;

    reg [15:0] mem[63:0];

    initial begin
        // // Teste 1: 35 + 50 - 62 + 50 = 72
        // mem[0] = 16'b1010000000100010; // LDI R0, 34
        // mem[1] = 16'b1010010000110010; // LDI R1, 50
        // mem[2] = 16'b0000000010000000; // ADD R0 = R0 + R1
        // mem[3] = 16'b1010100000111110; // LDI R2, 62
        // mem[4] = 16'b0010000100000000; // SUB R0 = R0 - R2
        // mem[5] = 16'b0000000010000000; // ADD R0 = R0 + R1
        // mem[6] = 16'b1110110000000000; // REP R3 = R0
        // mem[7] = 16'b1000110000000000; // OUT R3
        // mem[8] = 16'b0110000000000000; // HALT

        // Teste 2: 6 * 6 = 36
        mem[0] = 16'b1010010000000001; // LDI R1, 1
        mem[1] = 16'b1010100000000101; // LDI R2, 5
        mem[2] = 16'b1010110000000110; // LDI R3, 6
        mem[3] = 16'b1111000110000000; // REP R4 = R3
        mem[4] = 16'b0000111000000000; // ADD R3 = R3 + R4
        mem[5] = 16'b0010100010000000; // SUB R2 = R2 - R1
        mem[6] = 16'b1100100000000010; // BNE R2 2
        mem[7] = 16'b1100001111111101; // BNE R0 -3
        mem[8] = 16'b1000110000000000; // OUT R3
        mem[9] = 16'b0110000000000000; // HALT
    end

    always @(pc) begin
        out = mem[pc];
    end
endmodule